`ifdef tcm_defined

 `else 
`define tcm_defined
typedef int tcm;
`endif 
