
//************************************************************
//                                                            
//      Copyright Mentor Graphics Corporation 2006 - 2011     
//                  All Rights Reserved                       
//                                                            
//       THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY      
//         INFORMATION WHICH IS THE PROPERTY OF MENTOR        
//         GRAPHICS CORPORATION OR ITS LICENSORS AND IS       
//                 SUBJECT TO LICENSE TERMS.                  
//                                                            
//************************************************************


// Generated by Model Builder 

module ahb_slave_protocol
#(string	__portPath = "",
parameter	int	__portCount = 0,
parameter	string	__snapshotPath = "",
parameter	int	__timeFactor = 1
)

  (
    input DUMMY, 
    (*	master	*)	input	HSEL, 
    (*	master	*)	input	[1:0]	HTRANS	/* isAddress = 0 */, 
    (*	master	*)	input	HWRITE, 
    (*	master	*)	input	[63:0]	HADDR	/* isAddress = 1 */, 
    (*	master	=	2	*)	input	[2:0]	HSIZE	/* isAddress = 0 */, 
    (*	slave	=	0	*)	input	[1:0]	HRESP	/* isAddress = 0 */, 
    (*	slave	*)	input	[63:0]	HRDATA	/* isAddress = 0 */, 
    (*	master	*)	input	[63:0]	HWDATA	/* isAddress = 0 */, 
    (*	master	=	0	*)	input	[2:0]	HBURST	/* isAddress = 0 */, 
    (*	slave	*)	input	HREADY, 
    (*	clk	*)	input	CLK
  );

chandle __pMessageHandler;
chandle __pPort;
import "DPI-C" pure function void Papoulis_ReadVCD_ProtocolError(input string reason, input string functionName, input longint unsigned stime, input chandle pMessageHandler);

`ifdef OPEN_ARRAYS  
import "DPI-C" function void Papoulis_ReadVCD_SendMessage(
`else
import "DPI-C" function void Papoulis_ReadVCD_OldSendMessage(
`endif
input chandle pMessageHandler, input chandle pPort, input string messageName, input longint unsigned stime
`ifdef OPEN_ARRAYS  
, input longint unsigned paramArray []
`else
, input longint unsigned p1, input longint unsigned p2, input longint unsigned p3, input longint unsigned p4
`endif
);


import "DPI-C" function chandle Papoulis_ReadVCD_GetPortHandle(input chandle pMessageHandler, input string portPath);
import "DPI-C" function chandle Papoulis_ReadVCD_GetMessageHandler(input string snapshotPath, input int factor);


import "DPI-C" pure function int Papoulis_ReadVCD_CycleTimeSet(input chandle pMessageHandler, input string portPath, input longint unsigned low, input longint unsigned high);
import "DPI-C" pure function void Papoulis_ReadVCD_SaveCycleClkTime( input chandle pMessageHandler, input chandle pPort, input longint unsigned low, input longint unsigned high);
task findCycleTime();
    time currentTime;
    time lowTime;
    time highTime;
    integer isAlreadySet; 
    
    isAlreadySet	=	0;
begin
    while (!isAlreadySet) 
    begin
        @(negedge CLK);
        currentTime = $time;
        @(posedge CLK);
        lowTime = $time - currentTime;
        currentTime = $time;
        @(negedge CLK);
        highTime = $time - currentTime;
        isAlreadySet = Papoulis_ReadVCD_CycleTimeSet(__pMessageHandler, __portPath, lowTime, highTime);
    end
    Papoulis_ReadVCD_SaveCycleClkTime(__pMessageHandler, __pPort, lowTime, highTime);
end
endtask

initial
	findCycleTime();

typedef enum int {wait_nonseq_req=0, wait_write_ack, seq_write_or_end, 
wait_read_ack, write_data, end_sequence, seq_read_or_end}  PROTOCOL_STATES;

function void NONSEQ_WRITE_REQ(input longint unsigned HADDR, input longint unsigned HSIZE, input longint unsigned HBURST, input longint unsigned block_size);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = HADDR;
	paramArray[1] = HSIZE;
	paramArray[2] = HBURST;
	paramArray[3] = block_size;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "NONSEQ_WRITE_REQ", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "NONSEQ_WRITE_REQ", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, HADDR, HSIZE, HBURST, block_size
`endif
);
endfunction


function void WRITE_DATA(input longint unsigned HWDATA);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = HWDATA;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "WRITE_DATA", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "WRITE_DATA", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, HWDATA, 0, 0, 0
`endif
);
endfunction


function void SEQ_WRITE_REQ(input longint unsigned HADDR, input longint unsigned HSIZE, input longint unsigned block_size);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = HADDR;
	paramArray[1] = HSIZE;
	paramArray[2] = block_size;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "SEQ_WRITE_REQ", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "SEQ_WRITE_REQ", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, HADDR, HSIZE, block_size, 0
`endif
);
endfunction


function void NONSEQ_READ_REQ(input longint unsigned HADDR, input longint unsigned HSIZE, input longint unsigned HBURST, input longint unsigned block_size);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = HADDR;
	paramArray[1] = HSIZE;
	paramArray[2] = HBURST;
	paramArray[3] = block_size;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "NONSEQ_READ_REQ", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "NONSEQ_READ_REQ", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, HADDR, HSIZE, HBURST, block_size
`endif
);
endfunction


function void SEQ_READ_REQ(input longint unsigned HADDR, input longint unsigned HSIZE, input longint unsigned block_size);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = HADDR;
	paramArray[1] = HSIZE;
	paramArray[2] = block_size;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "SEQ_READ_REQ", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "SEQ_READ_REQ", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, HADDR, HSIZE, block_size, 0
`endif
);
endfunction


function void write_ack();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "write_ack", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "write_ack", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0
`endif
);
endfunction


function void bus_error();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "bus_error", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "bus_error", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0
`endif
);
endfunction


function void bus_split();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "bus_split", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "bus_split", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0
`endif
);
endfunction


function void bus_retry();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "bus_retry", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "bus_retry", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0
`endif
);
endfunction


function void END_TRANSACTION();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "END_TRANSACTION", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "END_TRANSACTION", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0
`endif
);
endfunction


function void read_ack(input longint unsigned HRDATA);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = HRDATA;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "read_ack", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "read_ack", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, HRDATA, 0, 0, 0
`endif
);
endfunction


function void protocolError;
input str;
string str;
$display(str);
Papoulis_ReadVCD_ProtocolError(str, "protocolError", $time, __pMessageHandler);
endfunction

PROTOCOL_STATES protocolState;
reg [2:0] HSIZE_reg;
int i;
always
    @(HSIZE)
        begin 
            HSIZE_reg = HSIZE;
            for(i = 0;(i<=2);i = (i + 1))
                begin 
                    if ((HSIZE_reg[i]===1'bz))
                    begin 
                        HSIZE_reg[i] = 1'b0;
                    end
                end
        end
(* protocol_initial *)
initial
    protocolState = wait_nonseq_req;
initial
begin
    __pMessageHandler = Papoulis_ReadVCD_GetMessageHandler(__snapshotPath, __timeFactor);
    __pPort = Papoulis_ReadVCD_GetPortHandle(__pMessageHandler, __portPath);
    while(1)
begin 
    case (protocolState)
    wait_nonseq_req:
        begin 
            if (((HSEL&&(HTRANS==2'b10))&&(HWRITE==1'b1)))
            begin 
                protocolState = write_data;
                (* WRITE *)
                NONSEQ_WRITE_REQ(HADDR,HSIZE_reg,HBURST,(1 << HSIZE_reg));
                @(negedge CLK)
                    ;
            end
            else
                if (((HSEL&&(HTRANS==2'b10))&&(HWRITE==1'b0)))
                begin 
                    protocolState = wait_read_ack;
                    (* READ *)
                    NONSEQ_READ_REQ(HADDR,HSIZE_reg,HBURST,(1 << HSIZE_reg));
                    @(negedge CLK)
                        ;
                end
                else
                    if ((HSEL!==1'b1))
                    begin 
                        protocolState = wait_nonseq_req;
                        @(negedge CLK)
                            ;
                    end
                    else
                        if ((HSEL&&(HTRANS==2'b00)))
                        begin 
                            protocolState = wait_nonseq_req;
                            @(negedge CLK)
                                ;
                        end
                        else
                        begin 
                            $display("protocol ahb_slave sequence is wrong, in state wait_nonseq_req\n");
                            $display("\tthere is no transition that possible at time: ",$time,"\n");
                            @(negedge CLK)
                                ;
                        end
        end
    write_data:
        begin 
            protocolState = wait_write_ack;
            WRITE_DATA(HWDATA);
        end
    wait_write_ack:
        begin 
            if ((!HREADY))
            begin 
                protocolState = wait_write_ack;
                @(negedge CLK)
                    ;
            end
            else
                if ((HRESP==2'b00))
                begin 
                    protocolState = seq_write_or_end;
                    write_ack();
                end
                else
                    if ((HRESP==2'b01))
                    begin 
                        protocolState = end_sequence;
                        bus_error();
                    end
                    else
                        if ((HRESP==2'b10))
                        begin 
                            protocolState = end_sequence;
                            bus_retry();
                        end
                        else
                            if ((HRESP==2'b11))
                            begin 
                                protocolState = end_sequence;
                                bus_split();
                            end
        end
    seq_write_or_end:
        begin 
            if ((HSEL&&(HTRANS==2'b01)))
            begin 
                protocolState = seq_write_or_end;
                @(negedge CLK)
                    ;
            end
            else
                if ((((HSEL&&(HTRANS==2'b10))||(HTRANS==2'b00))||(!HSEL)))
                begin 
                    protocolState = wait_nonseq_req;
                    END_TRANSACTION();
                end
                else
                begin 
                    protocolState = write_data;
                    SEQ_WRITE_REQ(HADDR,HSIZE_reg,(1 << HSIZE_reg));
                    @(negedge CLK)
                        ;
                end
        end
    wait_read_ack:
        begin 
            if ((!HREADY))
            begin 
                protocolState = wait_read_ack;
                @(negedge CLK)
                    ;
            end
            else
                if ((HRESP==2'b00))
                begin 
                    protocolState = seq_read_or_end;
                    read_ack(HRDATA);
                end
                else
                    if ((HRESP==2'b01))
                    begin 
                        protocolState = end_sequence;
                        bus_error();
                    end
                    else
                        if ((HRESP==2'b10))
                        begin 
                            protocolState = end_sequence;
                            bus_retry();
                        end
                        else
                            if ((HRESP==2'b11))
                            begin 
                                protocolState = end_sequence;
                                bus_split();
                            end
        end
    seq_read_or_end:
        begin 
            if ((HSEL&&(HTRANS==2'b01)))
            begin 
                protocolState = seq_read_or_end;
                @(negedge CLK)
                    ;
            end
            else
                if ((((HSEL&&(HTRANS==2'b10))||(HTRANS==2'b00))||(!HSEL)))
                begin 
                    protocolState = wait_nonseq_req;
                    END_TRANSACTION();
                end
                else
                begin 
                    protocolState = wait_read_ack;
                    SEQ_READ_REQ(HADDR,HSIZE_reg,(1 << HSIZE_reg));
                    @(negedge CLK)
                        ;
                end
        end
    end_sequence:
        begin 
            if ((((HSEL&&(HTRANS==2'b10))||(HTRANS==2'b00))||(!HSEL)))
            begin 
                protocolState = wait_nonseq_req;
                END_TRANSACTION();
            end
            else
            begin 
                $display("protocol ahb_slave sequence is wrong, in state end_read\n");
                $display("\tthere is no transition that possible at time: ",$time,"\n");
                @(negedge CLK)
                    ;
            end
        end
    endcase
end
end
endmodule
