`ifdef generic_defined

 `else 
`define generic_defined
typedef int generic;
`endif 
