
//************************************************************
//                                                            
//      Copyright Mentor Graphics Corporation 2006 - 2011     
//                  All Rights Reserved                       
//                                                            
//       THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY      
//         INFORMATION WHICH IS THE PROPERTY OF MENTOR        
//         GRAPHICS CORPORATION OR ITS LICENSORS AND IS       
//                 SUBJECT TO LICENSE TERMS.                  
//                                                            
//************************************************************


// Generated by Model Builder 

module axi_protocol
#(
    parameter WORD_SIZE = 32, 
    string	__portPath = "",
    parameter	int	__portCount = 0,
    parameter	string	__snapshotPath = "",
    parameter	int	__timeFactor = 1
)

  (
    input DUMMY, 
    (*	clk	*)	input	ACLK, 
    (*	master	*)	input	[3:0]	AWID	/* isAddress = 0 */, 
    (*	master	*)	input	[31:0]	AWADDR	/* isAddress = 1 */, 
    (*	master	*)	input	[3:0]	AWLEN	/* isAddress = 0 */, 
    (*	master	*)	input	[2:0]	AWSIZE	/* isAddress = 0 */, 
    (*	master	*)	input	[1:0]	AWBURST	/* isAddress = 0 */, 
    (*	master	*)	input	[1:0]	AWLOCK	/* isAddress = 0 */, 
    (*	master	*)	input	[3:0]	AWCACHE	/* isAddress = 0 */, 
    (*	master	*)	input	[2:0]	AWPROT	/* isAddress = 0 */, 
    (*	master	*)	input	AWVALID, 
    (*	slave	*)	input	AWREADY, 
    (*	master	*)	input	[3:0]	WID	/* isAddress = 0 */, 
    (*	master	*)	input	WLAST, 
    (*	master	*)	input	[WORD_SIZE - 1:0]	WDATA	/* isAddress = 0 */, 
    (*	master	*)	input	[WORD_SIZE / 8 - 1:0]	WSTRB	/* isAddress = 0 */, 
    (*	master	*)	input	WVALID, 
    (*	slave	*)	input	WREADY, 
    (*	slave	*)	input	[3:0]	BID	/* isAddress = 0 */, 
    (*	slave	*)	input	[1:0]	BRESP	/* isAddress = 0 */, 
    (*	slave	*)	input	BVALID, 
    (*	master	*)	input	BREADY, 
    (*	master	*)	input	[3:0]	ARID	/* isAddress = 0 */, 
    (*	master	*)	input	[31:0]	ARADDR	/* isAddress = 1 */, 
    (*	master	*)	input	[3:0]	ARLEN	/* isAddress = 0 */, 
    (*	master	*)	input	[2:0]	ARSIZE	/* isAddress = 0 */, 
    (*	master	*)	input	[1:0]	ARBURST	/* isAddress = 0 */, 
    (*	master	*)	input	[1:0]	ARLOCK	/* isAddress = 0 */, 
    (*	master	*)	input	[3:0]	ARCACHE	/* isAddress = 0 */, 
    (*	master	*)	input	[2:0]	ARPROT	/* isAddress = 0 */, 
    (*	master	*)	input	ARVALID, 
    (*	slave	*)	input	ARREADY, 
    (*	slave	*)	input	[3:0]	RID	/* isAddress = 0 */, 
    (*	slave	*)	input	RLAST, 
    (*	slave	*)	input	[WORD_SIZE - 1:0]	RDATA	/* isAddress = 0 */, 
    (*	slave	*)	input	[1:0]	RRESP	/* isAddress = 0 */, 
    (*	slave	*)	input	RVALID, 
    (*	master	*)	input	RREADY, 
    (*	master	*)	input	CACTIVE, 
    (*	slave	*)	input	CSYSREQ, 
    (*	master	*)	input	CSYSACK
  );

chandle __pMessageHandler;
chandle __pPort;
import "DPI-C" pure function void Papoulis_ReadVCD_ProtocolError(input string reason, input string functionName, input longint unsigned stime, input chandle pMessageHandler);

`ifdef OPEN_ARRAYS  
import "DPI-C" function void Papoulis_ReadVCD_SendMessage(
`else
import "DPI-C" function void Papoulis_ReadVCD_OldSendMessage(
`endif
input chandle pMessageHandler, input chandle pPort, input string messageName, input longint unsigned stime
`ifdef OPEN_ARRAYS  
, input longint unsigned paramArray []
`else
, input longint unsigned p1, input longint unsigned p2, input longint unsigned p3, input longint unsigned p4, input longint unsigned p5, input longint unsigned p6, input longint unsigned p7, input longint unsigned p8, input longint unsigned p9
`endif
);


import "DPI-C" function chandle Papoulis_ReadVCD_GetPortHandle(input chandle pMessageHandler, input string portPath);
import "DPI-C" function chandle Papoulis_ReadVCD_GetMessageHandler(input string snapshotPath, input int factor);


import "DPI-C" pure function int Papoulis_ReadVCD_CycleTimeSet(input chandle pMessageHandler, input string portPath, input longint unsigned low, input longint unsigned high);
import "DPI-C" pure function void Papoulis_ReadVCD_SaveCycleClkTime( input chandle pMessageHandler, input chandle pPort, input longint unsigned low, input longint unsigned high);
task findCycleTime();
    time currentTime;
    time lowTime;
    time highTime;
    integer isAlreadySet; 
    
    isAlreadySet	=	0;
begin
    while (!isAlreadySet) 
    begin
        @(negedge ACLK);
        currentTime = $time;
        @(posedge ACLK);
        lowTime = $time - currentTime;
        currentTime = $time;
        @(negedge ACLK);
        highTime = $time - currentTime;
        isAlreadySet = Papoulis_ReadVCD_CycleTimeSet(__pMessageHandler, __portPath, lowTime, highTime);
    end
    Papoulis_ReadVCD_SaveCycleClkTime(__pMessageHandler, __pPort, lowTime, highTime);
end
endtask

initial
	findCycleTime();


function void writeBurst_Control(input longint unsigned TR_ID, input longint unsigned AWADDR, input longint unsigned AWLEN, input longint unsigned AWSIZE, input longint unsigned block_size, input longint unsigned AWBURST, input longint unsigned AWLOCK, input longint unsigned AWCACHE, input longint unsigned AWPROT);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = TR_ID;
	paramArray[1] = AWADDR;
	paramArray[2] = AWLEN;
	paramArray[3] = AWSIZE;
	paramArray[4] = block_size;
	paramArray[5] = AWBURST;
	paramArray[6] = AWLOCK;
	paramArray[7] = AWCACHE;
	paramArray[8] = AWPROT;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "writeBurst_Control", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "writeBurst_Control", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, TR_ID, AWADDR, AWLEN, AWSIZE, block_size, AWBURST, AWLOCK, AWCACHE, AWPROT
`endif
);
$display($time," Master : Write Burst Control initiated ");
endfunction


function void writeBurst_Ready();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = 1;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "writeBurst_Ready", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "writeBurst_Ready", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 1, 0, 0, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Slave : Write Burst Control accepted ");
endfunction


function void writeBurst_Data(input longint unsigned TR_ID, input longint unsigned WDATA, input longint unsigned WSTRB);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = TR_ID;
	paramArray[1] = WDATA;
	paramArray[2] = WSTRB;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "writeBurst_Data", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "writeBurst_Data", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, TR_ID, WDATA, WSTRB, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Master : Write Burst Data initiated ");
endfunction


function void writeBurst_acceptData();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "writeBurst_acceptData", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "writeBurst_acceptData", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Slave : Write Burst Data accepted ");
endfunction


function void writeBurst_LastData(input longint unsigned TR_ID, input longint unsigned WDATA, input longint unsigned WSTRB);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = TR_ID;
	paramArray[1] = WDATA;
	paramArray[2] = WSTRB;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "writeBurst_LastData", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "writeBurst_LastData", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, TR_ID, WDATA, WSTRB, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Master : Write Burst Last Data initiated ");
endfunction


function void writeBurst_acceptLastData();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "writeBurst_acceptLastData", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "writeBurst_acceptLastData", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Slave : Write Burst Last Data accepted ");
endfunction


function void writeBurst_Response(input longint unsigned TR_ID, input longint unsigned BRESP);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = TR_ID;
	paramArray[1] = BRESP;
	paramArray[2] = 0;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "writeBurst_Response", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "writeBurst_Response", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, TR_ID, BRESP, 0, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Slave : Write Burst Response ");
endfunction


function void writeBurst_acceptResponse();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "writeBurst_acceptResponse", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "writeBurst_acceptResponse", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Master : Write Burst Response accepted ");
endfunction


function void writeBurst_Done();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "writeBurst_Done", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "writeBurst_Done", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Master : Write Burst Completed ");
endfunction


function void readBurst_Control(input longint unsigned TR_ID, input longint unsigned ARADDR, input longint unsigned ARLEN, input longint unsigned ARSIZE, input longint unsigned block_size, input longint unsigned ARBURST, input longint unsigned ARLOCK, input longint unsigned ARCACHE, input longint unsigned ARPROT);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = TR_ID;
	paramArray[1] = ARADDR;
	paramArray[2] = ARLEN;
	paramArray[3] = ARSIZE;
	paramArray[4] = block_size;
	paramArray[5] = ARBURST;
	paramArray[6] = ARLOCK;
	paramArray[7] = ARCACHE;
	paramArray[8] = ARPROT;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "readBurst_Control", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "readBurst_Control", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, TR_ID, ARADDR, ARLEN, ARSIZE, block_size, ARBURST, ARLOCK, ARCACHE, ARPROT
`endif
);
$display($time," Master : Read Burst Control initiated ");
endfunction


function void readBurst_Ready();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = 1;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "readBurst_Ready", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "readBurst_Ready", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 1, 0, 0, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Slave : Read Burst Control accepted ");
endfunction


function void readBurst_Data(input longint unsigned TR_ID, input longint unsigned RDATA, input longint unsigned RRESP);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = TR_ID;
	paramArray[1] = RDATA;
	paramArray[2] = RRESP;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "readBurst_Data", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "readBurst_Data", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, TR_ID, RDATA, RRESP, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Slave : Read Burst Data initiated ");
endfunction


function void readBurst_acceptData();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "readBurst_acceptData", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "readBurst_acceptData", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Master : Read Burst Data accepted ");
endfunction


function void readBurst_LastData(input longint unsigned TR_ID, input longint unsigned RDATA, input longint unsigned RRESP);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = TR_ID;
	paramArray[1] = RDATA;
	paramArray[2] = RRESP;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "readBurst_LastData", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "readBurst_LastData", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, TR_ID, RDATA, RRESP, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Slave : Read Burst Last Data initiated ");
endfunction


function void readBurst_acceptLastData();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "readBurst_acceptLastData", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "readBurst_acceptLastData", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Master : Read Burst Last Data accepted ");
endfunction


function void readBurst_Done();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 8];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
	paramArray[4] = 0;
	paramArray[5] = 0;
	paramArray[6] = 0;
	paramArray[7] = 0;
	paramArray[8] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "readBurst_Done", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "readBurst_Done", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0, 0, 0, 0, 0, 0
`endif
);
$display($time," Master : Read Burst Completed ");
endfunction

int ROutstanding = 0;
int WOutstanding = 0;
int WResponseOutstanding = 0;
logic [3:0] LockedID;
reg [3:0] WIDs[1:15] ;
reg AddrNeed[1:15] ;
int flag;
int i;
int j;
int RLockedAccessViolation_flag = 0;
int WLockedAccessViolation_flag = 0;
typedef enum int {UnLocked=0, Locked, LockLast}  LOCK_STATES;
LOCK_STATES LockState;
initial
    LockState = UnLocked;
typedef enum int {wait_writeAddress_req=0, wait_writeAddress_ack, 
wait_writeData_req, wait_writeData_ack, wait_writeLastData_ack, 
wait_loop_writeData_req, wait_writeResponse_req, wait_writeResponse_ack, 
end_write, wait_readAddress_req, wait_readAddress_ack, wait_readData_req, 
wait_readData_ack, wait_loop_readData_req, wait_readLastData_ack, end_read}  
PROTOCOL_STATES;
PROTOCOL_STATES AWprotocolState;
PROTOCOL_STATES WprotocolState;
PROTOCOL_STATES BprotocolState;
PROTOCOL_STATES ARprotocolState;
PROTOCOL_STATES RprotocolState;
(* SM_successor = wait_writeData_req *)
(* tlm_phase_start = "begin_req" *)
(* tlm_phase_end = "end_req" *)
(* protocol_initial *)
initial
    AWprotocolState = wait_writeAddress_req;
(* SM_successor = wait_writeResponse_req *)
(* protocol_initial *)
(* tlm_phase_start = "begin_resp" *)
(* tlm_phase_end = "end_resp" *)
initial
    WprotocolState = wait_writeData_req;
(* protocol_initial *)
initial
    BprotocolState = wait_writeResponse_req;
(* SM_successor = wait_readData_req *)
(* tlm_phase_start = "begin_req" *)
(* tlm_phase_end = "end_req" *)
(* protocol_initial *)
initial
    ARprotocolState = wait_readAddress_req;
(* protocol_initial *)
(* tlm_phase_start = "begin_resp" *)
(* tlm_phase_end = "end_resp" *)
initial
    RprotocolState = wait_readData_req;
always
    @(negedge ACLK)
        begin 
            if ((((AWVALID==1)&&(WLockedAccessViolation_flag==0))&&(AWREADY==1)))
            begin 
                if ((WOutstanding==0))
                begin 
                    WOutstanding++;
                    WIDs[WOutstanding] = AWID;
                end
                else
                begin 
                    flag = 0;
                    for(i = 1;(i<=WOutstanding);i = (i + 1))
                        begin 
                            if ((WIDs[i]==AWID))
                            begin 
                                flag = 1;
                                AddrNeed[i] = 0;
                            end
                        end
                    if ((flag==0))
                    begin 
                        WOutstanding++;
                        WIDs[WOutstanding] = AWID;
                    end
                end
            end
        end
always
    @(negedge ACLK)
        begin 
            if (((WVALID==1)&&(WREADY==1)))
            begin 
                if ((WOutstanding==0))
                begin 
                    WOutstanding++;
                    WIDs[WOutstanding] = WID;
                    AddrNeed[WOutstanding] = 1;
                end
                else
                begin 
                    flag = 0;
                    for(i = 1;(i<=WOutstanding);i = (i + 1))
                        begin 
                            if ((WIDs[i]==WID))
                            begin 
                                flag = 1;
                            end
                        end
                    if ((flag==0))
                    begin 
                        WOutstanding++;
                        WIDs[WOutstanding] = WID;
                        AddrNeed[WOutstanding] = 1;
                    end
                end
            end
        end
always
    @(negedge ACLK)
        begin 
            if (((BVALID==1)&&(BREADY==1)))
            begin 
                for(i = 1;(i<=WOutstanding);i = (i + 1))
                    begin 
                        if ((WIDs[i]==BID))
                            for(j = i;(j < WOutstanding);j = (j + 1))
                                begin 
                                    WIDs[j] = WIDs[(j + 1)];
                                    AddrNeed[j] = AddrNeed[(j + 1)];
                                end
                    end
            end
        end
always
    @(AWVALID)
        begin 
            if ((AWVALID===0))
                WLockedAccessViolation_flag = 0;
            else
                if ((AWVALID==1))
                begin 
                    case (LockState)
                    UnLocked:
                        if ((AWLOCK==2'b10))
                            if ((((ROutstanding==0)&&(WOutstanding==0))&&(~(((!$isunknown(ARVALID))&&
                            ARVALID)&&(ARLOCK!=2'b10)))))
                            begin 
                                LockState = Locked;
                                LockedID = AWID;
                                (* LockAccess *)
                                WLockedAccessViolation_flag = 0;
                            end
                            else
                            begin 
                                $display(
                                "Error: A master must wait for all outstanding transactions to complete before issuing a write address which is the first in a locked sequence."
                                );
                                WLockedAccessViolation_flag = 1;
                            end
                    Locked:
                        if ((AWID==LockedID))
                        begin 
                            if ((AWLOCK!=2'b10))
                                if ((((ROutstanding==0)&&(WOutstanding==0))&&(ARVALID!==1)))
                                begin 
                                    LockState = LockLast;
                                    (* UnLockAccess *)
                                    WLockedAccessViolation_flag = 0;
                                end
                                else
                                begin 
                                    $display(
                                    "Error: A master must wait for all locked transactions to complete before issuing an unlocked write address."
                                    );
                                    WLockedAccessViolation_flag = 1;
                                end
                        end
                        else
                        begin 
                            $display(
                            "Error: A master must ensure that all transactions within a locked sequence have the same ARID or AWID"
                            );
                            WLockedAccessViolation_flag = 1;
                        end
                    LockLast:
                        if ((((ROutstanding==0)&&(WOutstanding==0))&&(~((!$isunknown(ARVALID))&&(
                        ARVALID & (ARLOCK!=AWLOCK))))))
                        begin 
                            if ((AWLOCK==2'b10))
                            begin 
                                LockState = Locked;
                                LockedID = AWID;
                            end
                            else
                            begin 
                                LockState = UnLocked;
                                WLockedAccessViolation_flag = 0;
                            end
                        end
                        else
                        begin 
                            $display(
                            "Error: A master must wait for an unlocked transaction at the end of a locked sequence to complete before issuing another write address."
                            );
                            WLockedAccessViolation_flag = 1;
                        end
                    endcase
                end
        end
always
    @(ARVALID)
        begin 
            if ((ARVALID===0))
                RLockedAccessViolation_flag = 0;
            else
                if ((ARVALID===1))
                begin 
                    case (LockState)
                    UnLocked:
                        if ((ARLOCK==2'b10))
                            if ((((ROutstanding==0)&&(WOutstanding==0))&&(~(((!$isunknown(AWVALID))&&
                            AWVALID)&&(AWLOCK!=2'b10)))))
                            begin 
                                LockState = Locked;
                                LockedID = ARID;
                                (* LockAccess *)
                                RLockedAccessViolation_flag = 0;
                            end
                            else
                            begin 
                                $display(
                                "Error: A master must wait for all outstanding transactions to complete before issuing a read address which is the first in a locked sequence."
                                );
                                RLockedAccessViolation_flag = 1;
                            end
                    Locked:
                        if ((ARID==LockedID))
                        begin 
                            if ((ARLOCK!=2'b10))
                                if ((((ROutstanding==0)&&(WOutstanding==0))&&(AWVALID!==1)))
                                begin 
                                    LockState = LockLast;
                                    (* UnLockAccess *)
                                    RLockedAccessViolation_flag = 0;
                                end
                                else
                                begin 
                                    $display(
                                    "Error: A master must wait for all locked transactions to complete before issuing an unlocked read address."
                                    );
                                    RLockedAccessViolation_flag = 1;
                                end
                        end
                        else
                        begin 
                            $display(
                            "Error: A master must ensure that all transactions within a locked sequence have the same ARID or AWID"
                            );
                            RLockedAccessViolation_flag = 1;
                        end
                    LockLast:
                        if ((((ROutstanding==0)&&(WOutstanding==0))&&(~((!$isunknown(AWVALID))&&(
                        AWVALID & (AWLOCK!=ARLOCK))))))
                        begin 
                            if ((ARLOCK==2'b10))
                            begin 
                                LockState = Locked;
                                LockedID = ARID;
                            end
                            else
                            begin 
                                LockState = UnLocked;
                                RLockedAccessViolation_flag = 0;
                            end
                        end
                        else
                        begin 
                            $display(
                            "Error: A master must wait for an unlocked transaction at the end of a locked sequence to complete before issuing another read address."
                            );
                            RLockedAccessViolation_flag = 1;
                        end
                    endcase
                end
        end
initial
begin
    __pMessageHandler = Papoulis_ReadVCD_GetMessageHandler(__snapshotPath, __timeFactor);
    __pPort = Papoulis_ReadVCD_GetPortHandle(__pMessageHandler, __portPath);
    while(1)
begin 
    case (AWprotocolState)
    wait_writeAddress_req:
        begin 
            if (((AWVALID===1)&&(WLockedAccessViolation_flag==0)))
            begin 
                AWprotocolState = wait_writeAddress_ack;
                (* WRITE *)
                writeBurst_Control(AWID,AWADDR,AWLEN,AWSIZE,(1 << AWSIZE),AWBURST,AWLOCK,
                AWCACHE,AWPROT);
            end
            else
            begin 
                AWprotocolState = wait_writeAddress_req;
                @(negedge ACLK)
                    ;
            end
        end
    wait_writeAddress_ack:
        begin 
            if ((AWREADY===1))
            begin 
                AWprotocolState = wait_writeAddress_req;
                writeBurst_Ready();
                @(negedge ACLK)
                    ;
            end
            else
            begin 
                AWprotocolState = wait_writeAddress_ack;
                @(negedge ACLK)
                    ;
            end
        end
    endcase
end
end
initial
begin
    __pMessageHandler = Papoulis_ReadVCD_GetMessageHandler(__snapshotPath, __timeFactor);
    __pPort = Papoulis_ReadVCD_GetPortHandle(__pMessageHandler, __portPath);
    while(1)
begin 
    case (WprotocolState)
    wait_writeData_req:
        begin 
            if ((WVALID===1))
            begin 
                if ((WLAST===1))
                begin 
                    WprotocolState = wait_writeLastData_ack;
                    writeBurst_LastData(WID,WDATA,WSTRB);
                end
                else
                begin 
                    WprotocolState = wait_writeData_ack;
                    writeBurst_Data(WID,WDATA,WSTRB);
                end
            end
            else
            begin 
                WprotocolState = wait_writeData_req;
                @(negedge ACLK)
                    ;
            end
        end
    wait_loop_writeData_req:
        begin 
            if ((WVALID===1))
            begin 
                if ((WLAST===1))
                begin 
                    WprotocolState = wait_writeLastData_ack;
                    writeBurst_LastData(WID,WDATA,WSTRB);
                end
                else
                begin 
                    WprotocolState = wait_writeData_ack;
                    writeBurst_Data(WID,WDATA,WSTRB);
                end
            end
            else
            begin 
                WprotocolState = wait_loop_writeData_req;
                @(negedge ACLK)
                    ;
            end
        end
    wait_writeLastData_ack:
        begin 
            if ((WREADY===1))
            begin 
                WprotocolState = wait_writeData_req;
                writeBurst_acceptLastData();
                WResponseOutstanding++;
                @(negedge ACLK)
                    ;
            end
            else
            begin 
                WprotocolState = wait_writeLastData_ack;
                @(negedge ACLK)
                    ;
            end
        end
    wait_writeData_ack:
        begin 
            if ((WREADY===1))
            begin 
                if ((WLAST!==1))
                begin 
                    WprotocolState = wait_loop_writeData_req;
                    writeBurst_acceptData();
                    @(negedge ACLK)
                        ;
                end
            end
            else
            begin 
                WprotocolState = wait_writeData_ack;
                @(negedge ACLK)
                    ;
            end
        end
    endcase
end
end
initial
begin
    __pMessageHandler = Papoulis_ReadVCD_GetMessageHandler(__snapshotPath, __timeFactor);
    __pPort = Papoulis_ReadVCD_GetPortHandle(__pMessageHandler, __portPath);
    while(1)
begin 
    case (BprotocolState)
    wait_writeResponse_req:
        begin 
            if (((WResponseOutstanding!==0)&&(BVALID===1)))
            begin 
                BprotocolState = wait_writeResponse_ack;
                writeBurst_Response(BID,BRESP);
            end
            else
            begin 
                BprotocolState = wait_writeResponse_req;
                @(negedge ACLK)
                    ;
            end
        end
    wait_writeResponse_ack:
        begin 
            if ((BREADY===1))
            begin 
                BprotocolState = end_write;
                writeBurst_acceptResponse();
            end
            else
            begin 
                BprotocolState = wait_writeResponse_ack;
                @(negedge ACLK)
                    ;
            end
        end
    end_write:
        begin 
            BprotocolState = wait_writeResponse_req;
            writeBurst_Done();
            WResponseOutstanding--;
            WOutstanding--;
            @(negedge ACLK)
                ;
        end
    endcase
end
end
initial
begin
    __pMessageHandler = Papoulis_ReadVCD_GetMessageHandler(__snapshotPath, __timeFactor);
    __pPort = Papoulis_ReadVCD_GetPortHandle(__pMessageHandler, __portPath);
    while(1)
begin 
    case (ARprotocolState)
    wait_readAddress_req:
        begin 
            if (((ARVALID===1)&&(RLockedAccessViolation_flag==0)))
            begin 
                ARprotocolState = wait_readAddress_ack;
                (* READ *)
                readBurst_Control(ARID,ARADDR,ARLEN,ARSIZE,(1 << ARSIZE),ARBURST,ARLOCK,
                ARCACHE,ARPROT);
            end
            else
            begin 
                ARprotocolState = wait_readAddress_req;
                @(negedge ACLK)
                    ;
            end
        end
    wait_readAddress_ack:
        begin 
            if ((ARREADY===1))
            begin 
                ARprotocolState = wait_readAddress_req;
                readBurst_Ready();
                ROutstanding++;
                @(negedge ACLK)
                    ;
            end
            else
            begin 
                ARprotocolState = wait_readAddress_ack;
                @(negedge ACLK)
                    ;
            end
        end
    endcase
end
end
initial
begin
    __pMessageHandler = Papoulis_ReadVCD_GetMessageHandler(__snapshotPath, __timeFactor);
    __pPort = Papoulis_ReadVCD_GetPortHandle(__pMessageHandler, __portPath);
    while(1)
begin 
    case (RprotocolState)
    wait_readData_req:
        begin 
            if (((ROutstanding!==0)&&(RVALID===1)))
            begin 
                if ((RLAST===1))
                begin 
                    RprotocolState = wait_readLastData_ack;
                    readBurst_LastData(RID,RDATA,RRESP);
                end
                else
                begin 
                    RprotocolState = wait_readData_ack;
                    readBurst_Data(RID,RDATA,RRESP);
                end
            end
            else
            begin 
                RprotocolState = wait_readData_req;
                @(negedge ACLK)
                    ;
            end
        end
    wait_readLastData_ack:
        begin 
            if ((RREADY===1))
            begin 
                RprotocolState = end_read;
                readBurst_acceptLastData();
            end
            else
            begin 
                RprotocolState = wait_readLastData_ack;
                @(negedge ACLK)
                    ;
            end
        end
    wait_loop_readData_req:
        begin 
            if (((ROutstanding!==0)&&(RVALID===1)))
            begin 
                if ((RLAST===1))
                begin 
                    RprotocolState = wait_readLastData_ack;
                    readBurst_LastData(RID,RDATA,RRESP);
                end
                else
                begin 
                    RprotocolState = wait_readData_ack;
                    readBurst_Data(RID,RDATA,RRESP);
                end
            end
            else
            begin 
                RprotocolState = wait_loop_readData_req;
                @(negedge ACLK)
                    ;
            end
        end
    wait_readData_ack:
        begin 
            if ((RREADY===1))
            begin 
                if ((RLAST!==1))
                begin 
                    RprotocolState = wait_loop_readData_req;
                    readBurst_acceptData();
                    @(negedge ACLK)
                        ;
                end
            end
            else
            begin 
                RprotocolState = wait_readData_ack;
                @(negedge ACLK)
                    ;
            end
        end
    end_read:
        begin 
            RprotocolState = wait_readData_req;
            readBurst_Done();
            ROutstanding--;
            @(negedge ACLK)
                ;
        end
    endcase
end
end
endmodule
