
//************************************************************
//                                                            
//      Copyright Mentor Graphics Corporation 2006 - 2011     
//                  All Rights Reserved                       
//                                                            
//       THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY      
//         INFORMATION WHICH IS THE PROPERTY OF MENTOR        
//         GRAPHICS CORPORATION OR ITS LICENSORS AND IS       
//                 SUBJECT TO LICENSE TERMS.                  
//                                                            
//************************************************************


// Generated by Model Builder 

module usb_protocol
#(
    parameter endpoint_type_param = 0, 
    string	__portPath = "",
    parameter	int	__portCount = 0,
    parameter	string	__snapshotPath = "",
    parameter	int	__timeFactor = 1
)

  (
    input DUMMY, 
    (*	master	*)	input	[1:0]	LINESTATE	/* isAddress = 0 */, 
    (*	master	*)	input	[1:0]	XCVRSEL	/* isAddress = 0 */, 
    (*	master	*)	input	TERMSEL, 
    (*	master	*)	input	RXACTIVE, 
    (*	master	*)	input	RXVALID, 
    (*	master	*)	input	TXREADY, 
    (*	slave	*)	input	TXVALID, 
    (*	master	=	0	*)	input	[15:0]	XDATAIN	/* isAddress = 0 */, 
    (*	slave	*)	input	[15:0]	XDATAOUT	/* isAddress = 0 */, 
    (*	clk	*)	input	XCLK
  );

chandle __pMessageHandler;
chandle __pPort;
import "DPI-C" pure function void Papoulis_ReadVCD_ProtocolError(input string reason, input string functionName, input longint unsigned stime, input chandle pMessageHandler);

`ifdef OPEN_ARRAYS  
import "DPI-C" function void Papoulis_ReadVCD_SendMessage(
`else
import "DPI-C" function void Papoulis_ReadVCD_OldSendMessage(
`endif
input chandle pMessageHandler, input chandle pPort, input string messageName, input longint unsigned stime
`ifdef OPEN_ARRAYS  
, input longint unsigned paramArray []
`else
, input longint unsigned p1, input longint unsigned p2, input longint unsigned p3, input longint unsigned p4
`endif
);


import "DPI-C" function chandle Papoulis_ReadVCD_GetPortHandle(input chandle pMessageHandler, input string portPath);
import "DPI-C" function chandle Papoulis_ReadVCD_GetMessageHandler(input string snapshotPath, input int factor);


import "DPI-C" pure function int Papoulis_ReadVCD_CycleTimeSet(input chandle pMessageHandler, input string portPath, input longint unsigned low, input longint unsigned high);
import "DPI-C" pure function void Papoulis_ReadVCD_SaveCycleClkTime( input chandle pMessageHandler, input chandle pPort, input longint unsigned low, input longint unsigned high);
task findCycleTime();
    time currentTime;
    time lowTime;
    time highTime;
    integer isAlreadySet; 
    
    isAlreadySet	=	0;
begin
    while (!isAlreadySet) 
    begin
        @(negedge XCLK);
        currentTime = $time;
        @(posedge XCLK);
        lowTime = $time - currentTime;
        currentTime = $time;
        @(negedge XCLK);
        highTime = $time - currentTime;
        isAlreadySet = Papoulis_ReadVCD_CycleTimeSet(__pMessageHandler, __portPath, lowTime, highTime);
    end
    Papoulis_ReadVCD_SaveCycleClkTime(__pMessageHandler, __pPort, lowTime, highTime);
end
endtask

initial
	findCycleTime();

integer hSize = 0;
integer address = 0;
integer end_point = 0;
integer hs = 0;
integer fs = 0;
integer isMaster = 0;
typedef enum int {UNSET=0, HS, FS}  MODE;
MODE mode = UNSET;
integer endpoint_type = endpoint_type_param;

function void transmit_data(input longint unsigned XDATAOUT);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = XDATAOUT;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "transmit_data", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "transmit_data", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, XDATAOUT, 0, 0, 0
`endif
);
endfunction


function void transmit_data_packet(input longint unsigned XDATAOUT);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = XDATAOUT;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "transmit_data_packet", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "transmit_data_packet", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, XDATAOUT, 0, 0, 0
`endif
);
endfunction


function void transmit_handshake_packet(input longint unsigned XDATAOUT);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = XDATAOUT;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "transmit_handshake_packet", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "transmit_handshake_packet", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, XDATAOUT, 0, 0, 0
`endif
);
endfunction


function void end_trans_data(input longint unsigned hSize);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = hSize;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "end_trans_data", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "end_trans_data", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, hSize, 0, 0, 0
`endif
);
endfunction


function void no_handshake();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "no_handshake", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "no_handshake", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0
`endif
);
endfunction


function void continue_bulk();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "continue_bulk", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "continue_bulk", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0
`endif
);
endfunction


function void end_receive_data(input longint unsigned hSize);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = hSize;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "end_receive_data", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "end_receive_data", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, hSize, 0, 0, 0
`endif
);
endfunction


function void receive_data(input longint unsigned XDATAIN);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = XDATAIN;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "receive_data", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "receive_data", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, XDATAIN, 0, 0, 0
`endif
);
endfunction


function void receive_control_data(input longint unsigned end_point);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = end_point;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "receive_control_data", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "receive_control_data", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, end_point, 0, 0, 0
`endif
);
endfunction


function void receive_data_packet(input longint unsigned XDATAIN);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = XDATAIN;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "receive_data_packet", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "receive_data_packet", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, XDATAIN, 0, 0, 0
`endif
);
endfunction


function void receive_handshake_packet(input longint unsigned XDATAIN);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = XDATAIN;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "receive_handshake_packet", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "receive_handshake_packet", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, XDATAIN, 0, 0, 0
`endif
);
endfunction


function void master_no_handshake();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "master_no_handshake", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "master_no_handshake", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0
`endif
);
endfunction


function void invalid_packet();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "invalid_packet", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "invalid_packet", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0
`endif
);
endfunction


function void master_continue_bulk();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "master_continue_bulk", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "master_continue_bulk", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0, 0
`endif
);
endfunction


function void start_transaction(input longint unsigned address, input longint unsigned mode_p, input longint unsigned endpoint_type_p, input longint unsigned block_size);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = address;
	paramArray[1] = mode_p;
	paramArray[2] = endpoint_type_p;
	paramArray[3] = block_size;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "start_transaction", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "start_transaction", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, address, mode_p, endpoint_type_p, block_size
`endif
);
endfunction


function void receive_in_token_packet(input longint unsigned address, input longint unsigned mode_p, input longint unsigned endpoint_type_p);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = address;
	paramArray[1] = mode_p;
	paramArray[2] = endpoint_type_p;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "receive_in_token_packet", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "receive_in_token_packet", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, address, mode_p, endpoint_type_p, 0
`endif
);
endfunction


function void receive_out_token_packet(input longint unsigned address, input longint unsigned mode_p, input longint unsigned endpoint_type_p);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = address;
	paramArray[1] = mode_p;
	paramArray[2] = endpoint_type_p;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "receive_out_token_packet", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "receive_out_token_packet", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, address, mode_p, endpoint_type_p, 0
`endif
);
endfunction


function void receive_setup_token_packet(input longint unsigned address, input longint unsigned mode_p, input longint unsigned endpoint_type_p);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = address;
	paramArray[1] = mode_p;
	paramArray[2] = endpoint_type_p;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "receive_setup_token_packet", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "receive_setup_token_packet", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, address, mode_p, endpoint_type_p, 0
`endif
);
endfunction


function void receive_sof_token_packet(input longint unsigned address, input longint unsigned mode_p, input longint unsigned endpoint_type_p);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = address;
	paramArray[1] = mode_p;
	paramArray[2] = endpoint_type_p;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "receive_sof_token_packet", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "receive_sof_token_packet", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, address, mode_p, endpoint_type_p, 0
`endif
);
endfunction


function void receive_ping_packet(input longint unsigned address, input longint unsigned mode_p, input longint unsigned endpoint_type_p);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 3];
	paramArray[0] = address;
	paramArray[1] = mode_p;
	paramArray[2] = endpoint_type_p;
	paramArray[3] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "receive_ping_packet", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "receive_ping_packet", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, address, mode_p, endpoint_type_p, 0
`endif
);
endfunction


function void protocolError;
input error;
string error;
$display(error);
Papoulis_ReadVCD_ProtocolError(error, "protocolError", $time, __pMessageHandler);
endfunction

typedef enum int {idle_state=0, state_0, state_6, state_8, state_9, state_11, 
state_14, state_16, state_17, state_18, state_35, state_36, state_37}  
PROTOCOL_STATES;
PROTOCOL_STATES protocolState;
(* protocol_initial *)
initial
    protocolState = idle_state;
initial
begin
    __pMessageHandler = Papoulis_ReadVCD_GetMessageHandler(__snapshotPath, __timeFactor);
    __pPort = Papoulis_ReadVCD_GetPortHandle(__pMessageHandler, __portPath);
    while(1)
begin 
    case (protocolState)
    idle_state:
        begin 
            hs = ((XCVRSEL==0)&&(TERMSEL==0));
            fs = ((XCVRSEL==1)&&(TERMSEL==1));
            if (hs)
                mode = HS;
            if (fs)
                mode = FS;
            if (isMaster)
            begin 
                @(negedge XCLK)
                    ;
            end
            else
                if ((((RXACTIVE!==1)||(RXVALID!==1))||(((((XDATAIN[7:0] !=105)&&(XDATAIN[7:
                0] !=165))&&(XDATAIN[7:0] !=225))&&(XDATAIN[7:0] !=45))&&(XDATAIN[7:0] !=180))))
                begin 
                    if ((TXVALID&&TXREADY))
                    begin 
                        protocolError(
                        "ERROR: The current usb protocol is for an usb slave, only a master can transmit from idle state"
                        );
                        isMaster = 1;
                        @(negedge XCLK)
                            ;
                    end
                    else
                    begin 
                        protocolState = idle_state;
                        @(negedge XCLK)
                            ;
                    end
                end
                else
                    if ((((((XDATAIN[7:0] ==105)||(XDATAIN[7:0] ==225))||(XDATAIN[7:0] ==45))||
                    (XDATAIN[7:0] ==165))||(XDATAIN[7:0] ==180)))
                    begin 
                        protocolState = state_0;
                        end_point = XDATAIN[15:15] ;
                        address = XDATAIN[14:8] ;
                        (* IN_PACKET *)
                        (* OUT_PACKET *)
                        (* SETUP_PACKET *)
                        (* SOF_PACKET *)
                        (* PING_PACKET *)
                        start_transaction(address,mode,endpoint_type,2);
                    end
                    else
                    begin 
                        protocolError(
                        "ERROR:\tprotocol usb sequence is wrong, in state idle_state\n\tthere is no transition that possible"
                        );
                        @(negedge XCLK)
                            ;
                    end
        end
    state_0:
        begin 
            end_point = XDATAIN[15:15] ;
            address = XDATAIN[14:8] ;
            if ((XDATAIN[7:0] ==105))
            begin 
                protocolState = state_6;
                (* IN_PACKET *)
                receive_in_token_packet(address,mode,endpoint_type);
                @(negedge XCLK)
                    ;
            end
            else
                if ((XDATAIN[7:0] ==225))
                begin 
                    protocolState = state_14;
                    (* OUT_PACKET *)
                    receive_out_token_packet(address,mode,endpoint_type);
                    @(negedge XCLK)
                        ;
                end
                else
                    if ((XDATAIN[7:0] ==45))
                    begin 
                        protocolState = state_14;
                        (* SETUP_PACKET *)
                        receive_setup_token_packet(address,mode,endpoint_type);
                        @(negedge XCLK)
                            ;
                    end
                    else
                        if ((XDATAIN[7:0] ==165))
                        begin 
                            protocolState = state_35;
                            (* SOF_PACKET *)
                            receive_sof_token_packet(address,mode,endpoint_type);
                            @(negedge XCLK)
                                ;
                        end
                        else
                            if ((XDATAIN[7:0] ==180))
                            begin 
                                protocolState = state_36;
                                (* PING_PACKET *)
                                receive_ping_packet(address,mode,endpoint_type);
                                @(negedge XCLK)
                                    ;
                            end
        end
    state_6:
        begin 
            if ((!RXVALID))
            begin 
                protocolState = state_6;
                @(negedge XCLK)
                    ;
            end
            else
                if (RXVALID)
                begin 
                    protocolState = state_8;
                    end_point = ((XDATAIN[2:0]  << 1) + end_point);
                    receive_control_data(end_point);
                    @(negedge XCLK)
                        ;
                end
                else
                begin 
                    protocolError(
                    "ERROR:\tprotocol usb sequence is wrong, in state state_6\n\tthere is no transition that possible"
                    );
                    @(negedge XCLK)
                        ;
                end
        end
    state_8:
        begin 
            if (((TXVALID===0)&&(RXACTIVE===0)))
            begin 
                protocolState = state_8;
                @(negedge XCLK)
                    ;
            end
            else
                if (RXACTIVE)
                begin 
                    protocolState = idle_state;
                    no_handshake();
                end
                else
                    if (TXVALID)
                    begin 
                        @(negedge XCLK)
                            ;
                        if (((((XDATAOUT[7:0] ==15)||(XDATAOUT[7:0] ==135))||(XDATAOUT[7:0] ==75))||(
                        XDATAOUT[7:0] ==195)))
                        begin 
                            protocolState = state_9;
                            transmit_data_packet(XDATAOUT);
                            @(negedge XCLK)
                                ;
                        end
                        else
                            if ((((XDATAOUT[7:0] ==90)||(XDATAOUT[7:0] ==30))||(XDATAOUT[7:0] ==150)))
                            begin 
                                protocolState = idle_state;
                                transmit_handshake_packet(XDATAOUT);
                                @(negedge XCLK)
                                    ;
                            end
                    end
                    else
                    begin 
                        protocolError(
                        "ERROR:\tprotocol usb sequence is wrong, in state state_8\n\tthere is no transition that possible"
                        );
                        @(negedge XCLK)
                            ;
                    end
        end
    state_9:
        begin 
            if ((!TXVALID))
            begin 
                protocolState = state_11;
                hSize = (XDATAOUT[7:0] ==XDATAOUT[15:8] );
                end_trans_data(hSize);
                @(negedge XCLK)
                    ;
            end
            else
                if ((!TXREADY))
                begin 
                    protocolState = state_9;
                    @(negedge XCLK)
                        ;
                end
                else
                begin 
                    protocolState = state_9;
                    transmit_data(XDATAOUT);
                    @(negedge XCLK)
                        ;
                end
        end
    state_11:
        begin 
            if ((endpoint_type==1))
            begin 
                protocolState = idle_state;
                master_no_handshake();
            end
            else
                if (((!RXVALID)||(!RXACTIVE)))
                begin 
                    protocolState = state_11;
                    @(negedge XCLK)
                        ;
                end
                else
                    if ((RXVALID&&((((XDATAIN[7:0] ==210)||(XDATAIN[7:0] ==90))||(XDATAIN[7:0] 
                    ==30))||(XDATAIN[7:0] ==150))))
                    begin 
                        protocolState = idle_state;
                        receive_handshake_packet(XDATAIN);
                        @(negedge XCLK)
                            ;
                    end
                    else
                        if (((endpoint_type==2)&&((XDATAIN[7:0] ==105)||(XDATAIN[7:0] ==225))))
                        begin 
                            protocolState = idle_state;
                            master_continue_bulk();
                        end
                        else
                        begin 
                            protocolError(
                            "protocol usb sequence is wrong, in state state_11\n\tthere is no transition that possible"
                            );
                            @(negedge XCLK)
                                ;
                        end
        end
    state_14:
        begin 
            if ((!RXVALID))
            begin 
                protocolState = state_14;
                @(negedge XCLK)
                    ;
            end
            else
                if (RXVALID)
                begin 
                    protocolState = state_16;
                    end_point = ((XDATAIN[2:0]  << 1) + end_point);
                    receive_control_data(end_point);
                    @(negedge XCLK)
                        ;
                end
                else
                begin 
                    protocolError(
                    "protocol usb sequence is wrong, in state state_14\n\tthere is no transition that possible"
                    );
                    @(negedge XCLK)
                        ;
                end
        end
    state_16:
        begin 
            if (((!RXACTIVE)||(!RXVALID)))
            begin 
                protocolState = state_16;
                @(negedge XCLK)
                    ;
            end
            else
                if ((RXVALID&&((((XDATAIN[7:0] ==195)||(XDATAIN[7:0] ==75))||(XDATAIN[7:0] 
                ==135))||(XDATAIN[7:0] ==15))))
                begin 
                    protocolState = state_17;
                    receive_data_packet(XDATAIN);
                    @(negedge XCLK)
                        ;
                end
                else
                begin 
                    protocolState = idle_state;
                    invalid_packet();
                end
        end
    state_17:
        begin 
            if (RXVALID)
            begin 
                protocolState = state_17;
                receive_data(XDATAIN);
                @(negedge XCLK)
                    ;
            end
            else
                if (((!RXACTIVE)&&((hs&&(LINESTATE[1:0] ==0))||(fs&&(LINESTATE[1:0] ==1)))))
                begin 
                    protocolState = state_18;
                    hSize = (XDATAIN[7:0] ==XDATAIN[15:8] );
                    end_receive_data(hSize);
                end
                else
                begin 
                    protocolState = state_17;
                    @(negedge XCLK)
                        ;
                end
        end
    state_18:
        begin 
            if ((endpoint_type==1))
            begin 
                protocolState = idle_state;
                no_handshake();
            end
            else
                if (((TXVALID===0)&&(RXACTIVE===0)))
                begin 
                    protocolState = state_18;
                    @(negedge XCLK)
                        ;
                end
                else
                    if (TXVALID)
                    begin 
                        @(negedge XCLK)
                            ;
                        if (((((XDATAOUT[7:0] ==210)||(XDATAOUT[7:0] ==90))||(XDATAOUT[7:0] ==30))||(
                        XDATAOUT[7:0] ==150)))
                        begin 
                            protocolState = idle_state;
                            transmit_handshake_packet(XDATAOUT);
                            @(negedge XCLK)
                                ;
                        end
                    end
                    else
                        if ((!RXVALID))
                        begin 
                            protocolState = state_18;
                            @(negedge XCLK)
                                ;
                        end
                        else
                            if (((endpoint_type==2)&&((XDATAIN[7:0] ==225)||(XDATAIN[7:0] ==105))))
                            begin 
                                protocolState = idle_state;
                                continue_bulk();
                            end
                            else
                            begin 
                                protocolError(
                                "protocol usb sequence is wrong, in state state_18\n\tthere is no transition that possible"
                                );
                                @(negedge XCLK)
                                    ;
                            end
        end
    state_35:
        begin 
            if ((!RXVALID))
            begin 
                protocolState = state_35;
                @(negedge XCLK)
                    ;
            end
            else
            begin 
                protocolState = idle_state;
                end_point = ((XDATAIN[2:0]  << 1) + end_point);
                receive_control_data(end_point);
            end
        end
    state_36:
        begin 
            if ((!RXVALID))
            begin 
                protocolState = state_36;
                @(negedge XCLK)
                    ;
            end
            else
                if (RXVALID)
                begin 
                    protocolState = state_37;
                    end_point = ((XDATAIN[2:0]  << 1) + end_point);
                    receive_control_data(end_point);
                    @(negedge XCLK)
                        ;
                end
                else
                begin 
                    protocolError(
                    "protocol usb sequence is wrong, in state state_14\n\tthere is no transition that possible"
                    );
                    @(negedge XCLK)
                        ;
                end
        end
    state_37:
        begin 
            if (RXACTIVE)
            begin 
                protocolState = idle_state;
                no_handshake();
            end
            else
                if (((TXVALID===0)&&(RXACTIVE===0)))
                begin 
                    protocolState = state_37;
                    @(negedge XCLK)
                        ;
                end
                else
                    if (TXVALID)
                    begin 
                        @(negedge XCLK)
                            ;
                        if (((((XDATAOUT[7:0] ==210)||(XDATAOUT[7:0] ==90))||(XDATAOUT[7:0] ==30))||(
                        XDATAOUT[7:0] ==150)))
                        begin 
                            protocolState = idle_state;
                            transmit_handshake_packet(XDATAOUT);
                            @(negedge XCLK)
                                ;
                        end
                    end
                    else
                    begin 
                        protocolError(
                        "protocol usb sequence is wrong, in state state_37\n\tthere is no transition that possible"
                        );
                        @(negedge XCLK)
                            ;
                    end
        end
    endcase
end
end
endmodule
