`ifdef usb_defined

 `else 
`define usb_defined
typedef int usb;
`endif 
