`ifdef ram_defined

 `else 
`define ram_defined
typedef int ram;
`endif 
