`ifdef axi_defined

 `else 
`define axi_defined
typedef int axi;
`endif 
