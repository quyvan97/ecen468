`ifdef ahb_master_defined

 `else 
`define ahb_master_defined
typedef int ahb_master;
`endif 
