`ifdef apb_defined

 `else 
`define apb_defined
typedef int apb;
`endif 
