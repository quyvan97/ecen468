`ifdef ahb_slave_defined

 `else 
`define ahb_slave_defined
typedef int ahb_slave;
`endif 
