
//************************************************************
//                                                            
//      Copyright Mentor Graphics Corporation 2006 - 2011     
//                  All Rights Reserved                       
//                                                            
//       THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY      
//         INFORMATION WHICH IS THE PROPERTY OF MENTOR        
//         GRAPHICS CORPORATION OR ITS LICENSORS AND IS       
//                 SUBJECT TO LICENSE TERMS.                  
//                                                            
//************************************************************


// Generated by Model Builder 

module ram_protocol
#(
    parameter ADDR_WIDTH = 19,
    parameter DATA_WIDTH = 8, 
    string	__portPath = "",
    parameter	int	__portCount = 0,
    parameter	string	__snapshotPath = "",
    parameter	int	__timeFactor = 1
)

  (
    input DUMMY, 
    (*	clk	*)	input	clk, 
    (*	master	*)	input	ram_we, 
    (*	master	*)	input	[ADDR_WIDTH - 1:0]	ram_addr	/* isAddress = 1 */, 
    (*	master	=	0	*)	input	[DATA_WIDTH - 1:0]	ram_data_in	/* isAddress = 0 */, 
    (*	slave	=	0	*)	input	[DATA_WIDTH - 1:0]	ram_data_out	/* isAddress = 0 */
  );

chandle __pMessageHandler;
chandle __pPort;
import "DPI-C" pure function void Papoulis_ReadVCD_ProtocolError(input string reason, input string functionName, input longint unsigned stime, input chandle pMessageHandler);

`ifdef OPEN_ARRAYS  
import "DPI-C" function void Papoulis_ReadVCD_SendMessage(
`else
import "DPI-C" function void Papoulis_ReadVCD_OldSendMessage(
`endif
input chandle pMessageHandler, input chandle pPort, input string messageName, input longint unsigned stime
`ifdef OPEN_ARRAYS  
, input longint unsigned paramArray []
`else
, input longint unsigned p1, input longint unsigned p2, input longint unsigned p3
`endif
);


import "DPI-C" function chandle Papoulis_ReadVCD_GetPortHandle(input chandle pMessageHandler, input string portPath);
import "DPI-C" function chandle Papoulis_ReadVCD_GetMessageHandler(input string snapshotPath, input int factor);


import "DPI-C" pure function int Papoulis_ReadVCD_CycleTimeSet(input chandle pMessageHandler, input string portPath, input longint unsigned low, input longint unsigned high);
import "DPI-C" pure function void Papoulis_ReadVCD_SaveCycleClkTime( input chandle pMessageHandler, input chandle pPort, input longint unsigned low, input longint unsigned high);
task findCycleTime();
    time currentTime;
    time lowTime;
    time highTime;
    integer isAlreadySet; 
    
    isAlreadySet	=	0;
begin
    while (!isAlreadySet) 
    begin
        @(negedge clk);
        currentTime = $time;
        @(posedge clk);
        lowTime = $time - currentTime;
        currentTime = $time;
        @(negedge clk);
        highTime = $time - currentTime;
        isAlreadySet = Papoulis_ReadVCD_CycleTimeSet(__pMessageHandler, __portPath, lowTime, highTime);
    end
    Papoulis_ReadVCD_SaveCycleClkTime(__pMessageHandler, __pPort, lowTime, highTime);
end
endtask

initial
	findCycleTime();


function void NONSEQ_WRITE(input longint unsigned ram_addr, input longint unsigned ram_data_in, input longint unsigned block_size);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 2];
	paramArray[0] = ram_addr;
	paramArray[1] = ram_data_in;
	paramArray[2] = block_size;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "NONSEQ_WRITE", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "NONSEQ_WRITE", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, ram_addr, ram_data_in, block_size
`endif
);
$display("%0t/I, %m :- NONSEQ_WRITE(ram_addr=%0h, ram_data_in=%0h)",$time,
ram_addr,ram_data_in);
endfunction


function void SEQ_WRITE(input longint unsigned ram_addr, input longint unsigned ram_data_in, input longint unsigned block_size);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 2];
	paramArray[0] = ram_addr;
	paramArray[1] = ram_data_in;
	paramArray[2] = block_size;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "SEQ_WRITE", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "SEQ_WRITE", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, ram_addr, ram_data_in, block_size
`endif
);
$display("%0t/I, %m :- SEQ_WRITE(ram_addr=%0h, ram_data_in=%0h)",$time,
ram_addr,ram_data_in);
endfunction


function void nonseq_write_ack();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 2];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "nonseq_write_ack", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "nonseq_write_ack", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0
`endif
);
$display("%0t/O, %m :- nonseq_write_ack()",$time);
endfunction


function void seq_write_ack(input longint unsigned addr_count);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 2];
	paramArray[0] = addr_count;
	paramArray[1] = 0;
	paramArray[2] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "seq_write_ack", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "seq_write_ack", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, addr_count, 0, 0
`endif
);
$display("%0t/O, %m :- seq_write_ack(addr_count=%0h)",$time,addr_count);
endfunction


function void NONSEQ_READ(input longint unsigned ram_addr, input longint unsigned block_size);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 2];
	paramArray[0] = ram_addr;
	paramArray[1] = block_size;
	paramArray[2] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "NONSEQ_READ", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "NONSEQ_READ", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, ram_addr, block_size, 0
`endif
);
$display("%0t/I, %m :- NONSEQ_READ(ram_addr=%0h)",$time,ram_addr);
endfunction


function void SEQ_READ(input longint unsigned ram_addr, input longint unsigned block_size);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 2];
	paramArray[0] = ram_addr;
	paramArray[1] = block_size;
	paramArray[2] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "SEQ_READ", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "SEQ_READ", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, ram_addr, block_size, 0
`endif
);
$display("%0t/I, %m :- SEQ_READ(ram_addr=%0h)",$time,ram_addr);
endfunction


function void nonseq_read_ack(input longint unsigned ram_data_out);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 2];
	paramArray[0] = ram_data_out;
	paramArray[1] = 0;
	paramArray[2] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "nonseq_read_ack", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "nonseq_read_ack", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, ram_data_out, 0, 0
`endif
);
$display("%0t/O, %m :- nonseq_read_ack(ram_data_out=%0h)",$time,ram_data_out);
endfunction


function void seq_read_ack(input longint unsigned ram_data_out, input longint unsigned addr_count);
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 2];
	paramArray[0] = ram_data_out;
	paramArray[1] = addr_count;
	paramArray[2] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "seq_read_ack", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "seq_read_ack", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, ram_data_out, addr_count, 0
`endif
);
$display("%0t/O, %m :- seq_read_ack(ram_data_out=%0h, addr_count=%0h)",$time,
ram_data_out,addr_count);
endfunction


function void END_TRANSACTION();
`ifdef OPEN_ARRAYS  
	longint unsigned paramArray [0 : 2];
	paramArray[0] = 0;
	paramArray[1] = 0;
	paramArray[2] = 0;
`endif
`ifdef OPEN_ARRAYS  
	Papoulis_ReadVCD_SendMessage(__pMessageHandler, __pPort, "END_TRANSACTION", $time
`else
	Papoulis_ReadVCD_OldSendMessage(__pMessageHandler, __pPort, "END_TRANSACTION", $time
`endif
`ifdef OPEN_ARRAYS  
, paramArray
`else
, 0, 0, 0
`endif
);
$display("%0t/I, %m :- END_TRANSACTION()",$time);
endfunction


function void protocolError;
input error;
string error;
$display($time," --> ERROR in %m");
Papoulis_ReadVCD_ProtocolError(error, "protocolError", $time, __pMessageHandler);
endfunction

reg [(ADDR_WIDTH - 1):0] start_ram_addr;
reg [(ADDR_WIDTH - 1):0] addr_count;
typedef enum int {IDLE=0, NONSEQ_WRITE_STATE, WRITE_LOOP_STATE, 
SEQ_WRITE_STATE, NONSEQ_READ_STATE, READ_LOOP_STATE, SEQ_READ_STATE}  
PROTOCOL_STATES;
PROTOCOL_STATES protocolState;
(* protocol_initial *)
initial
    protocolState = IDLE;
initial
begin
    __pMessageHandler = Papoulis_ReadVCD_GetMessageHandler(__snapshotPath, __timeFactor);
    __pPort = Papoulis_ReadVCD_GetPortHandle(__pMessageHandler, __portPath);
    while(1)
begin 
    case (protocolState)
    IDLE:
        begin 
            if (((((| ram_addr)===1'b0)||((| ram_addr)===1'bX))||((| ram_addr)===1'bZ)))
            begin 
                protocolState = IDLE;
                @(negedge clk)
                    ;
            end
            else
                if ((ram_we==1'b1))
                begin 
                    protocolState = NONSEQ_WRITE_STATE;
                    start_ram_addr = ram_addr;
                    (* WRITE *)
                    NONSEQ_WRITE(ram_addr,ram_data_in,1);
                    @(negedge clk)
                        ;
                end
                else
                    if ((ram_we==1'b0))
                    begin 
                        protocolState = NONSEQ_READ_STATE;
                        start_ram_addr = ram_addr;
                        (* READ *)
                        NONSEQ_READ(ram_addr,1);
                        @(negedge clk)
                            ;
                    end
                    else
                    begin 
                        protocolError("protocol ram sequence is wrong in state IDLE");
                        @(negedge clk)
                            ;
                    end
        end
    NONSEQ_WRITE_STATE:
        begin 
            protocolState = WRITE_LOOP_STATE;
            addr_count = 1'b0;
            nonseq_write_ack();
            @(negedge clk)
                ;
        end
    WRITE_LOOP_STATE:
        begin 
            if (((((| ram_addr)===1'b0)||((| ram_addr)===1'bX))||((| ram_addr)===1'bZ)))
            begin 
                protocolState = WRITE_LOOP_STATE;
                @(negedge clk)
                    ;
            end
            else
                if ((ram_addr==((start_ram_addr + addr_count) + 1'b1)))
                begin 
                    protocolState = SEQ_WRITE_STATE;
                    SEQ_WRITE(ram_addr,ram_data_in,1);
                    @(negedge clk)
                        ;
                end
                else
                begin 
                    protocolState = IDLE;
                    END_TRANSACTION();
                end
        end
    SEQ_WRITE_STATE:
        begin 
            protocolState = WRITE_LOOP_STATE;
            addr_count = (addr_count + 1'b1);
            seq_write_ack(addr_count);
            @(negedge clk)
                ;
        end
    NONSEQ_READ_STATE:
        begin 
            protocolState = READ_LOOP_STATE;
            addr_count = 1'b0;
            nonseq_read_ack(ram_data_out);
            @(negedge clk)
                ;
        end
    READ_LOOP_STATE:
        begin 
            if (((((| ram_addr)===1'b0)||((| ram_addr)===1'bX))||((| ram_addr)===1'bZ)))
            begin 
                protocolState = READ_LOOP_STATE;
                @(negedge clk)
                    ;
            end
            else
                if ((ram_addr==((start_ram_addr + addr_count) + 1'b1)))
                begin 
                    protocolState = SEQ_READ_STATE;
                    SEQ_READ(ram_addr,1);
                    @(negedge clk)
                        ;
                end
                else
                begin 
                    protocolState = IDLE;
                    END_TRANSACTION();
                end
        end
    SEQ_READ_STATE:
        begin 
            protocolState = READ_LOOP_STATE;
            addr_count = (addr_count + 1'b1);
            seq_read_ack(ram_data_out,addr_count);
            @(negedge clk)
                ;
        end
    endcase
end
end
endmodule
