`ifdef signal_defined

 `else 
`define signal_defined
typedef int signal;
`endif 
